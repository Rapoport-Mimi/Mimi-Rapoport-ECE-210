/*
 * Copyright (c) 2024 Mimi Rapoport
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_Rapoport (
    input  reg  [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out[6:0] = 0;
  assign uio_oe = 0;
  assign uo_out = 0;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, clk, rst_n, 1'b0};

  // Instantiate perceptron
  perceptron perceptron1 (
    .clk(clk), 
    .reset(rst_n), 
    .in1(ui_in[3:0]), 
    .in2(ui_in[7:4]), 
    .in3(uio_in[6:0]), 
    .desired_out(uio_in[7]), 
    .out(uio_out[7])
  );

endmodule
